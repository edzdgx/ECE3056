-- Edward Zhou / 903130547
-- control unit. simply implements the truth table for a small set of
-- instructions
--
-- added seT pc_Hazard value

Library IEEE;
use IEEE.std_logic_1164.all;

entity control is
port(opcode, ex_opcode: in std_logic_vector(5 downto 0);
     ex_wreg_addr : in std_logic_vector(4 downto 0);
     instruction : in std_logic_vector(31 downto 0);
     RegDst, MemRead, MemToReg, MemWrite, PC_HAZARD :out  std_logic;
     ALUSrc, RegWrite, Branch: out std_logic;
     ALUOp: out std_logic_vector(1 downto 0));
end control;

architecture behavioral of control is

signal rformat, lw, sw, beq  :std_logic; -- define local signals
				    -- corresponding to instruction
				    -- type

 begin
--
-- recognize opcode for each instruction type
-- these variable should be inferred as wires

	rformat     <=  '1'  WHEN  Opcode = "000000"  ELSE '0';
	Lw          <=  '1'  WHEN  Opcode = "100011"  ELSE '0';
 	Sw          <=  '1'  WHEN  Opcode = "101011"  ELSE '0';
   	Beq         <=  '1'  WHEN  Opcode = "000100"  ELSE '0';

-- if load && detection = '1'
PC_HAZARD <= '1' when (opcode ="000000" and ex_opcode = "100011" and ((ex_wreg_addr = instruction(25 downto 21) or ex_wreg_addr = instruction(20 downto 16)))) else '0';

--
-- implement each output signal as the column of the truth
-- table  which defines the control
--

RegDst <= rformat;
ALUSrc <= (lw or sw) ;

MemToReg <= lw ;
RegWrite <= (rformat or lw);
MemRead <= lw ;
MemWrite <= sw;
Branch <= beq;

ALUOp(1 downto 0) <=  rformat & '0'; -- note the use of the concatenation operator
				     -- to form  2 bit signal

end behavioral;
